LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
USE IEEE.STD_LOGIC_SIGNED.ALL;

ENTITY Adder IS
	PORT (
					input_0, input_1 : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
					output : OUT STD_LOGIC_VECTOR(15 DOWNTO 0)
				);
END ENTITY;

ARCHITECTURE behavioral OF Adder IS
BEGIN
	output <= input_0 + input_1;
END ARCHITECTURE;


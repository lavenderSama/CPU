LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
USE IEEE.STD_LOGIC_SIGNED.ALL;

ENTITY Pause IS
    PORT ( MEM      : IN STD_LOGIC_VECTOR(1 downto 0);
           LAST_TO_WRITE: IN STD_LOGIC_VECTOR(2 downto 0);
           NEXT10_8 : IN STD_LOGIC_VECTOR(2 downto 0);
           NEXT7_5  : IN STD_LOGIC_VECTOR(2 downto 0);
           NEXT15_0 : IN STD_LOGIC_VECTOR(15 downto 0);
           PAUSE_SIGNAL: OUT STD_LOGIC);
END Pause;

ARCHITECTURE behavior of Pause IS
BEGIN
	process (MEM, LAST_TO_WRITE, NEXT10_8, NEXT7_5, NEXT15_0)
	begin
    case MEM is
        when "10" => if (LAST_TO_WRITE = NEXT10_8) then
                        case NEXT15_0(15 downto 11) is
                            when "01001" => PAUSE_SIGNAL <='1'; --ADDIU
                            when "01000" => PAUSE_SIGNAL <='1'; --ADDIU3
                            when "11100" => PAUSE_SIGNAL <='1'; --ADDU,SUBU
                            when "11101" => case NEXT15_0(4 downto 0) is --AND,CMP,JR,MFPC,OR,JRRA,JALR
                                                 when "01100" | "01010" | "01101" => PAUSE_SIGNAL <='1';
                                                 when "00000" => --JR, MFPC, JRRA, JALR
                                                 	case NEXT15_0(7 downto 5) is
                                                 		when "000" | "110" => PAUSE_SIGNAL <= '1'; --JR, JALR
                                                 		when "001" | "010" => PAUSE_SIGNAL <= '0'; --JRRA, MFPC
                                                 		when others => PAUSE_SIGNAL <= '0';
                                                 	end case;
                                                 when "01011" => PAUSE_SIGNAL <= '0'; --NEG
                                                 when others => PAUSE_SIGNAL <='0';
                                            end case;
                            when "00100" => PAUSE_SIGNAL <='1'; --BEQZ
                            when "00101" => PAUSE_SIGNAL <='1'; --BNEZ
                            when "11110" =>  --MFIH,MTIH
                            	case NEXT15_0(0) is
								                when '0' =>  --MFIH
								                    PAUSE_SIGNAL <= '0';
								                when '1' =>  --MTIH
								                    PAUSE_SIGNAL <='1';
								                when others => PAUSE_SIGNAL <= '0';
								              end case;								                    
                            when "10011" => PAUSE_SIGNAL <='1'; --LW
                            when "11011" | "11010" => PAUSE_SIGNAL <='1'; --SW, SW_SP
                            when others => PAUSE_SIGNAL <='0';
                        end case;
                    elsif (LAST_TO_WRITE = NEXT7_5) then
                        case NEXT15_0(15 downto 11) is
                            when "11100" => PAUSE_SIGNAL <= '1'; --ADDU,SUBU
                            when "11101" => case NEXT15_0(4 downto 0) is --AND,CMP,JR,MFPC,OR,JRRA,JALR, NEG
                                              when "01100" | "01010" | "01101" | "01011" => PAUSE_SIGNAL <='1';
                                              when "00000" => --JR, MFPC, JRRA, JALR
                                               	PAUSE_SIGNAL <= '0';
                                              when others  => PAUSE_SIGNAL <='0';
                                            end case;
                            when "01111" => PAUSE_SIGNAL <= '1'; --MOVE
                            when "00110" => PAUSE_SIGNAL <= '1'; --SLL,SRA
                            when "01100" => if (NEXT15_0(10 downto 8) = "100") then --MTSP
                            									PAUSE_SIGNAL <= '1';
                            								else
                            									PAUSE_SIGNAL <= '0';
                            								end if;
                            when "11011" => PAUSE_SIGNAL <= '1';
                            when others => PAUSE_SIGNAL <='0';
                        end case;
                    else
                        PAUSE_SIGNAL<='0';
                    end if;
        when "00"|"01"|"11" => PAUSE_SIGNAL<='0';
		  when others => PAUSE_SIGNAL<='0';
    end case;
	end process;
END behavior;
